module defaults

pub const session_ttl = 60
