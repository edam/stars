module main

fn main() {
	mut app := App.new()
	app.run()
}
